module lab7_2(
   input clk,
   input rst,
   output [3:0] vgaRed,
   output [3:0] vgaGreen,
   output [3:0] vgaBlue,
   output hsync,
   output vsync,
    input up,
    input down,
    input left,
    input right,
    input hint,
    output reg pass
    );

integer i;
integer j;
integer k;

/*reg [0:63] init_cells = {
    4'd0,  4'd1,  4'd2,  4'd3,
    4'd4,  4'd5,  4'd6, 4'd7,
    4'd8, 4'd9,  4'd10, 4'd11,
    4'd12, 4'd13, 4'd14, 4'd15
};*/
reg [0:63] pass_cells = {
    4'd1,  4'd2,  4'd3,  4'd4,
    4'd5,  4'd6,  4'd7, 4'd8,
    4'd9, 4'd10,  4'd11, 4'd12,
    4'd13, 4'd14, 4'd15, 4'd0
};
reg [0:63] init_cells = {
    4'd2,  4'd3,  4'd4,  4'd8,
    4'd1,  4'd6,  4'd7, 4'd12,
    4'd5, 4'd10,  4'd0, 4'd11,
    4'd9, 4'd13, 4'd14, 4'd15
};

reg [0:63] cells ;
reg [0:63] next_cells;

parameter INIT = 2'd0;
parameter GAME = 2'd1;
parameter HINT = 2'd2;
parameter PASS = 2'd3;
reg [1:0] state = INIT;
reg [1:0] next_state;

reg next_pass;

wire clk_25MHz;
wire valid;
wire [9:0] h_cnt; //640
wire [9:0] v_cnt; //480

wire rst_debounced;
wire up_debounced;
wire down_debounced;
wire left_debounced;
wire right_debounced;

wire rst_1pulse;
wire up_1pulse;
wire down_1pulse;
wire left_1pulse;
wire right_1pulse;

my_debounce db1 (.pb_debounced(rst_debounced), .pb(rst), .clk(clk));
my_debounce db2 (.pb_debounced(up_debounced), .pb(up), .clk(clk));
my_debounce db3 (.pb_debounced(down_debounced), .pb(down), .clk(clk));
my_debounce db4 (.pb_debounced(left_debounced), .pb(left), .clk(clk));
my_debounce db5 (.pb_debounced(right_debounced), .pb(right), .clk(clk));

my_OnePulse op1 (.signal_single_pulse(rst_1pulse), .signal(rst_debounced), .clock(clk));
my_OnePulse op2 (.signal_single_pulse(up_1pulse), .signal(up_debounced), .clock(clk));
my_OnePulse op3 (.signal_single_pulse(down_1pulse), .signal(down_debounced), .clock(clk));
my_OnePulse op4 (.signal_single_pulse(left_1pulse), .signal(left_debounced), .clock(clk));
my_OnePulse op5 (.signal_single_pulse(right_1pulse), .signal(right_debounced), .clock(clk));

     clock_divider clk_wiz_0_inst(
      .clk(clk),
      .clk1(clk_25MHz)
    );

   my_pixel_gen pixel_gen_inst(
       .h_cnt(h_cnt),
       .valid(valid),
       .vgaRed(vgaRed),
       .vgaGreen(vgaGreen),
       .vgaBlue(vgaBlue),
       .v_cnt(v_cnt),
       .cells(hint == 1'b1 ? pass_cells : cells)
    );

    my_vga_controller   vga_inst(
      .pclk(clk_25MHz),
      .reset(rst_1pulse),
      .hsync(hsync),
      .vsync(vsync),
      .valid(valid),
      .h_cnt(h_cnt),
      .v_cnt(v_cnt)
    );
// STATE    
always @(posedge clk or posedge rst_1pulse) begin
    if(rst_1pulse) begin
        state <= INIT;
    end
    else begin
        state <= next_state;
    end
end

always @* begin
    next_state = state;
    case(state)
        INIT : begin
            next_state = GAME;
        end
        GAME : begin
            if(hint == 1'b1) begin
                next_state = HINT;
            end
            else if(pass == 1'b1) begin
                next_state = PASS;
            end
        end
        HINT : begin
            if(hint == 1'b0) begin
                next_state = GAME;
            end
        end
    endcase
end
// CELLS
always @(posedge clk or posedge rst_1pulse) begin
    if(rst_1pulse) begin
        cells <= init_cells;
    end
    else begin
        cells <= next_cells;
    end
end

always @* begin
    next_cells = cells;
    case(state)
        INIT : begin
            next_cells = init_cells;
        end
        GAME : begin
            if(up_1pulse) begin
                for(i=0; i<16; i=i+1) begin
                    if(cells[i*4 +: 4] == 4'd0) begin
                        j = i;
                    end
                end
                if(j >= 0 && j <= 11) begin
                    //j = i+4;
                    next_cells[(j+4)*4 +: 4] = 4'd0;
                    next_cells[j*4 +: 4] = cells[(j+4)*4 +: 4];
                end
            end
            else if(down_1pulse) begin
                for(i=0; i<16; i=i+1) begin
                    if(cells[i*4 +: 4] == 4'd0) begin
                        j = i;
                    end
                end
                if(j >= 4 && j <= 15) begin
                    //j = i-4;
                    next_cells[(j-4)*4 +: 4] = 4'd0;
                    next_cells[j*4 +: 4] = cells[(j-4)*4 +: 4];
                end
            end
            else if(left_1pulse) begin
                for(i=0; i<16; i=i+1) begin
                    if(cells[i*4 +: 4] == 4'd0) begin
                        j = i;
                    end
                end
                if(j%4 != 3) begin
                    //j = i+1;
                    next_cells[(j+1)*4 +: 4] = 4'd0;
                    next_cells[j*4 +: 4] = cells[(j+1)*4 +: 4];
                end
            end
            else if(right_1pulse) begin
                for(i=0; i<16; i=i+1) begin
                    if(cells[i*4 +: 4] == 4'd0) begin
                        j = i;
                    end
                end
                if(j%4 != 0) begin
                    //j = i-1;
                    next_cells[(j-1)*4 +: 4] = 4'd0;
                    next_cells[j*4 +: 4] = cells[(j-1)*4 +: 4];
                end
            end
        end
    endcase
end     
// PASS
always @(posedge clk or posedge rst_1pulse) begin
    if(rst_1pulse) begin
        pass <= 1'b0;
    end
    else begin
        pass <= next_pass;
    end
end

always @* begin
    next_pass = pass;
    case(state)
        INIT : begin
            next_pass = 1'b0;
        end
        GAME : begin
            next_pass = 1'b1;
            for(k=0; k<16; k=k+1) begin
                if(cells[k*4 +: 4] != pass_cells[k*4 +: 4]) begin
                    next_pass = 1'b0;
                end
            end
        end
    endcase
end
endmodule

module my_debounce (
	input wire clk,
	input wire pb, 
	output wire pb_debounced 
);
	reg [3:0] shift_reg; 

	always @(posedge clk) begin
		shift_reg[3:1] <= shift_reg[2:0];
		shift_reg[0] <= pb;
	end

	assign pb_debounced = ((shift_reg == 4'b1111) ? 1'b1 : 1'b0);

endmodule

module my_OnePulse (
	output reg signal_single_pulse,
	input wire signal,
	input wire clock
	);
	
	reg signal_delay;

	always @(posedge clock) begin
		if (signal == 1'b1 & signal_delay == 1'b0)
		  signal_single_pulse <= 1'b1;
		else
		  signal_single_pulse <= 1'b0;

		signal_delay <= signal;
	end
endmodule

module my_pixel_gen(
   input [9:0] h_cnt,
   input valid,
   output reg [3:0] vgaRed,
   output reg [3:0] vgaGreen,
   output reg [3:0] vgaBlue,
   input [9:0] v_cnt,
   input [0:63] cells
   );

// div 8, >> 3
// 640 -> 80 / 4 = 20
// 480 -> 60 / 4 = 15

parameter [11:0] position [0:15] = {
    12'd0, 12'd20, 12'd40, 12'd60,
    12'd1200, 12'd1220, 12'd1240, 12'd1260,
    12'd2400, 12'd2420, 12'd2440, 12'd2460,
    12'd3600, 12'd3620, 12'd3640, 12'd3660
};

parameter [11:0] color [0:4799] = {
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'hFFF,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000,
12'h000
};
     
always @(*) begin
    if(!valid)
        {vgaRed, vgaGreen, vgaBlue} = 12'h0;
    else if(v_cnt < 120) begin
        if(h_cnt < 160)
            {vgaRed, vgaGreen, vgaBlue} = color[position[cells[0:3]] + ((v_cnt>>3)%15)*80 + (h_cnt>>3)%20];
        else if(h_cnt < 320)
            {vgaRed, vgaGreen, vgaBlue} = color[position[cells[4:7]] + ((v_cnt>>3)%15)*80 + (h_cnt>>3)%20];
        else if(h_cnt < 480)
            {vgaRed, vgaGreen, vgaBlue} = color[position[cells[8:11]] + ((v_cnt>>3)%15)*80 + (h_cnt>>3)%20];
        else if(h_cnt < 640)
            {vgaRed, vgaGreen, vgaBlue} = color[position[cells[12:15]] + ((v_cnt>>3)%15)*80 + (h_cnt>>3)%20];
        else
            {vgaRed, vgaGreen, vgaBlue} = 12'h000;
    end
    else if(v_cnt < 240) begin
        if(h_cnt < 160)
            {vgaRed, vgaGreen, vgaBlue} = color[position[cells[16:19]] + ((v_cnt>>3)%15)*80 + (h_cnt>>3)%20];
        else if(h_cnt < 320)
            {vgaRed, vgaGreen, vgaBlue} = color[position[cells[20:23]] + ((v_cnt>>3)%15)*80 + (h_cnt>>3)%20];
        else if(h_cnt < 480)
            {vgaRed, vgaGreen, vgaBlue} = color[position[cells[24:27]] + ((v_cnt>>3)%15)*80 + (h_cnt>>3)%20];
        else if(h_cnt < 640)
            {vgaRed, vgaGreen, vgaBlue} = color[position[cells[28:31]] + ((v_cnt>>3)%15)*80 + (h_cnt>>3)%20];
        else
            {vgaRed, vgaGreen, vgaBlue} = 12'h000;
    end
    else if(v_cnt < 360) begin
        if(h_cnt < 160)
            {vgaRed, vgaGreen, vgaBlue} = color[position[cells[32:35]] + ((v_cnt>>3)%15)*80 + (h_cnt>>3)%20];
        else if(h_cnt < 320)
            {vgaRed, vgaGreen, vgaBlue} = color[position[cells[36:39]] + ((v_cnt>>3)%15)*80 + (h_cnt>>3)%20];
        else if(h_cnt < 480)
            {vgaRed, vgaGreen, vgaBlue} = color[position[cells[40:43]] + ((v_cnt>>3)%15)*80 + (h_cnt>>3)%20];
        else if(h_cnt < 640)
            {vgaRed, vgaGreen, vgaBlue} = color[position[cells[44:47]] + ((v_cnt>>3)%15)*80 + (h_cnt>>3)%20];
        else
            {vgaRed, vgaGreen, vgaBlue} = 12'h000;
    end
    else if(v_cnt < 480) begin
        if(h_cnt < 160)
            {vgaRed, vgaGreen, vgaBlue} = color[position[cells[48:51]] + ((v_cnt>>3)%15)*80 + (h_cnt>>3)%20];
        else if(h_cnt < 320)
            {vgaRed, vgaGreen, vgaBlue} = color[position[cells[52:55]] + ((v_cnt>>3)%15)*80 + (h_cnt>>3)%20];
        else if(h_cnt < 480)
            {vgaRed, vgaGreen, vgaBlue} = color[position[cells[56:59]] + ((v_cnt>>3)%15)*80 + (h_cnt>>3)%20];
        else if(h_cnt < 640)
            {vgaRed, vgaGreen, vgaBlue} = color[position[cells[60:63]] + ((v_cnt>>3)%15)*80 + (h_cnt>>3)%20];
        else
            {vgaRed, vgaGreen, vgaBlue} = 12'h000;
    end
    else
         {vgaRed, vgaGreen, vgaBlue} = 12'h0;
end
endmodule

`timescale 1ns/1ps
/////////////////////////////////////////////////////////////////
// Module Name: vga
/////////////////////////////////////////////////////////////////

module my_vga_controller (
    input wire pclk, reset,
    output wire hsync, vsync, valid,
    output wire [9:0]h_cnt,
    output wire [9:0]v_cnt
    );

    reg [9:0]pixel_cnt;
    reg [9:0]line_cnt;
    reg hsync_i,vsync_i;

    parameter HD = 640;
    parameter HF = 16;
    parameter HS = 96;
    parameter HB = 48;
    parameter HT = 800; 
    parameter VD = 480;
    parameter VF = 10;
    parameter VS = 2;
    parameter VB = 33;
    parameter VT = 525;
    parameter hsync_default = 1'b1;
    parameter vsync_default = 1'b1;

    always @(posedge pclk)
        if (reset)
            pixel_cnt <= 0;
        else
            if (pixel_cnt < (HT - 1))
                pixel_cnt <= pixel_cnt + 1;
            else
                pixel_cnt <= 0;

    always @(posedge pclk)
        if (reset)
            hsync_i <= hsync_default;
        else
            if ((pixel_cnt >= (HD + HF - 1)) && (pixel_cnt < (HD + HF + HS - 1)))
                hsync_i <= ~hsync_default;
            else
                hsync_i <= hsync_default; 

    always @(posedge pclk)
        if (reset)
            line_cnt <= 0;
        else
            if (pixel_cnt == (HT -1))
                if (line_cnt < (VT - 1))
                    line_cnt <= line_cnt + 1;
                else
                    line_cnt <= 0;

    always @(posedge pclk)
        if (reset)
            vsync_i <= vsync_default; 
        else if ((line_cnt >= (VD + VF - 1)) && (line_cnt < (VD + VF + VS - 1)))
            vsync_i <= ~vsync_default; 
        else
            vsync_i <= vsync_default; 

    assign hsync = hsync_i;
    assign vsync = vsync_i;
    assign valid = ((pixel_cnt < HD) && (line_cnt < VD));

    assign h_cnt = (pixel_cnt < HD) ? pixel_cnt : 10'd0;
    assign v_cnt = (line_cnt < VD) ? line_cnt : 10'd0;

endmodule
